  module encoder_256_8 (
    input  logic [239:0] interrupt_accepted,
    output logic [7:0]   sel_enc  
);

    logic            [255:0] temp_256   ;  
    localparam logic [7:0]   BASE = 8'd0;

    assign temp_256 = {16'b0,interrupt_accepted};

  always_comb begin 
    case (temp_256)
     // 256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + ;
      
      // Output for reserved from 253 to 158
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001: sel_enc = BASE + 0     ; // 255 - 255 

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002: sel_enc = BASE + 2-1   ; // 255 - 255 + 1

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004: sel_enc = BASE + 3-1   ; //253

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0008: sel_enc = BASE + 4-1   ; //252
      
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010: sel_enc = BASE + 5-1   ; //251

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0020: sel_enc = BASE + 6-1   ; //250

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0040: sel_enc = BASE + 7-1   ; //249
  
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0080: sel_enc = BASE + 8-1   ; //248
     
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100: sel_enc = BASE + 9-1   ; //247

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0200: sel_enc = BASE + 10-1  ; //246

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0400: sel_enc = BASE + 11-1  ; //245

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0800: sel_enc = BASE + 12-1  ; //244
      
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000: sel_enc = BASE + 13-1  ; //243

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_2000: sel_enc = BASE + 14-1  ; //242

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000: sel_enc = BASE + 15-1  ; //241

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_8000: sel_enc = BASE + 16-1  ; //240

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000: sel_enc = BASE + 17-1  ; //239

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000: sel_enc = BASE + 18-1  ; //238

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000: sel_enc = BASE + 19-1  ; //237

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0008_0000: sel_enc = BASE + 20-1  ; //236

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000: sel_enc = BASE + 21-1  ; //235

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0020_0000: sel_enc = BASE + 22-1  ; //234

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0040_0000: sel_enc = BASE + 23-1  ; //233

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0080_0000: sel_enc = BASE + 24-1  ; //232
 
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000: sel_enc = BASE + 25-1  ; //231

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0200_0000: sel_enc = BASE + 26-1  ; //230

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0400_0000: sel_enc = BASE + 27-1  ; //229

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000: sel_enc = BASE + 28-1  ; //228
     
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000: sel_enc = BASE + 29-1  ; //227

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_2000_0000: sel_enc = BASE + 30-1  ; //226

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0000: sel_enc = BASE + 31-1  ; //225

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_8000_0000: sel_enc = BASE + 32-1  ; //224
     
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000: sel_enc = BASE + 33-1  ; //223

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000: sel_enc = BASE + 34-1  ; //222

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000: sel_enc = BASE + 35-1  ; //221

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0008_0000_0000: sel_enc = BASE + 36-1  ; //220

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000: sel_enc = BASE + 37-1  ; //219

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0020_0000_0000: sel_enc = BASE + 38-1  ; //218

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0040_0000_0000: sel_enc = BASE + 39-1  ; //217

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0080_0000_0000: sel_enc = BASE + 40-1  ; //216
    
      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000: sel_enc = BASE + 41-1  ; //215

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0200_0000_0000: sel_enc = BASE + 42-1  ; //214

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0400_0000_0000: sel_enc = BASE + 43-1  ; //213

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0000: sel_enc = BASE + 44-1  ; //212

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000: sel_enc = BASE + 45-1  ; //211

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_2000_0000_0000: sel_enc = BASE + 46-1  ; //210

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0000_0000: sel_enc = BASE + 47-1  ; //209

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_8000_0000_0000: sel_enc = BASE + 48-1  ; //208

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000: sel_enc = BASE + 49-1  ; //207

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000: sel_enc = BASE + 50-1  ; //206

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000: sel_enc = BASE + 51-1  ; //205

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0008_0000_0000_0000: sel_enc = BASE + 52-1  ; //204

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000: sel_enc = BASE + 53-1  ; //203

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0020_0000_0000_0000: sel_enc = BASE + 54-1  ; //202

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0040_0000_0000_0000: sel_enc = BASE + 55-1  ; //201

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0080_0000_0000_0000: sel_enc = BASE + 56-1  ; //200

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000: sel_enc = BASE + 57-1  ; //199

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0200_0000_0000_0000: sel_enc = BASE + 58-1  ; //198

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0400_0000_0000_0000: sel_enc = BASE + 59-1  ; //197

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0000_0000: sel_enc = BASE + 60-1  ; //196

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000: sel_enc = BASE + 61-1  ; //195

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_2000_0000_0000_0000: sel_enc = BASE + 62-1  ; //194

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0000_0000_0000: sel_enc = BASE + 63-1  ; //193

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_8000_0000_0000_0000: sel_enc = BASE + 64-1  ; //192

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000: sel_enc = BASE + 65-1  ; //191

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000: sel_enc = BASE + 66-1  ; //190

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000: sel_enc = BASE + 67-1  ; //189

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0008_0000_0000_0000_0000: sel_enc = BASE + 68-1  ; //188

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000: sel_enc = BASE + 69-1  ; //187

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0020_0000_0000_0000_0000: sel_enc = BASE + 70-1  ; //186

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0040_0000_0000_0000_0000: sel_enc = BASE + 71-1  ; //185

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0080_0000_0000_0000_0000: sel_enc = BASE + 72-1  ; //184

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000: sel_enc = BASE + 73-1  ; //183

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0200_0000_0000_0000_0000: sel_enc = BASE + 74-1  ; //182

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0400_0000_0000_0000_0000: sel_enc = BASE + 75-1  ; //181

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0000_0000_0000: sel_enc = BASE + 76-1  ; //180

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000: sel_enc = BASE + 77-1  ; //179

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_2000_0000_0000_0000_0000: sel_enc = BASE + 78-1  ; //178

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000: sel_enc = BASE + 79-1  ; //177

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_8000_0000_0000_0000_0000: sel_enc = BASE + 80-1  ; //176

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000: sel_enc = BASE + 81-1  ; //175

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000: sel_enc = BASE + 82-1  ; //174

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000: sel_enc = BASE + 83-1  ; //173

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0008_0000_0000_0000_0000_0000: sel_enc = BASE + 84-1  ; //172

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000: sel_enc = BASE + 85-1  ; //171

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0020_0000_0000_0000_0000_0000: sel_enc = BASE + 86-1  ; //170

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0040_0000_0000_0000_0000_0000: sel_enc = BASE + 87-1  ; //169

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0080_0000_0000_0000_0000_0000: sel_enc = BASE + 88-1  ; //168

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000: sel_enc = BASE + 89-1  ; //167

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000: sel_enc = BASE + 90-1  ; //166

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0400_0000_0000_0000_0000_0000: sel_enc = BASE + 91-1  ; //165

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0000_0000_0000_0000: sel_enc = BASE + 92-1  ; //164

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000: sel_enc = BASE + 93-1  ; //163

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_2000_0000_0000_0000_0000_0000: sel_enc = BASE + 94-1  ; //162

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000: sel_enc = BASE + 95-1  ; //161

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_8000_0000_0000_0000_0000_0000: sel_enc = BASE + 96-1  ; //160

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 97-1  ;  //159

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 98-1  ; //158

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 99-1  ; //157

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0008_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 100-1 ; //156

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 101-1 ; //155

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0020_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 102-1 ; //154

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0040_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 103-1 ; //153

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0080_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 104-1 ; //152

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 105-1 ; //151

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 106-1 ; //150

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0400_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 107-1 ; //149

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 108-1 ; //148

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 109-1 ; //147

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_2000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 110-1 ; //146

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 111-1 ; //145

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0000_8000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 112-1 ; //144

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 113-1 ; //143

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 114-1 ; //142

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 115-1 ; //141

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0008_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 116-1 ; //140

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 117-1 ; //139

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0020_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 118-1 ; //138

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0040_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 119-1 ; //137

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0080_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 120-1 ; //136

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 121-1 ; //135

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 122-1 ; //134

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0400_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 123-1 ; //133

      256'h0000_0000_0000_0000_0000_0000_0000_0000_0800_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 124-1 ; //132

      256'h0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 125-1 ; //131

      256'h0000_0000_0000_0000_0000_0000_0000_0000_2000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 126-1 ; //130

      256'h0000_0000_0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 127-1 ; //129

      256'h0000_0000_0000_0000_0000_0000_0000_0000_8000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 128-1 ; //128

      256'h0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 129-1 ; //127

      256'h0000_0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 130-1 ; //126

      256'h0000_0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 131-1 ; //125

      256'h0000_0000_0000_0000_0000_0000_0000_0008_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 132-1 ; //124

      256'h0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 133-1 ; //123

      256'h0000_0000_0000_0000_0000_0000_0000_0020_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 134-1 ; //122

      256'h0000_0000_0000_0000_0000_0000_0000_0040_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 135-1 ; //121

      256'h0000_0000_0000_0000_0000_0000_0000_0080_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 136-1 ; //120

      256'h0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 137-1 ; //119

      256'h0000_0000_0000_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 138-1 ; //118

      256'h0000_0000_0000_0000_0000_0000_0000_0400_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 139-1 ; //117

      256'h0000_0000_0000_0000_0000_0000_0000_0800_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 140-1 ; //116

      256'h0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 141-1 ; //115

      256'h0000_0000_0000_0000_0000_0000_0000_2000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 142-1 ; //114

      256'h0000_0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 143-1 ; //113

      256'h0000_0000_0000_0000_0000_0000_0000_8000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 144-1 ; //112

      256'h0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 145-1 ; //111

      256'h0000_0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 146-1 ; //110

      256'h0000_0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 147-1 ; //109

      256'h0000_0000_0000_0000_0000_0000_0008_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 148-1 ; //108

      256'h0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 149-1 ; //107

      256'h0000_0000_0000_0000_0000_0000_0020_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 150-1 ; //106

      256'h0000_0000_0000_0000_0000_0000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 151-1 ; //105

      256'h0000_0000_0000_0000_0000_0000_0080_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 152-1 ; //104

      256'h0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 153-1 ; //103

      256'h0000_0000_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 154-1 ; //102

      256'h0000_0000_0000_0000_0000_0000_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 155-1 ; //101

      256'h0000_0000_0000_0000_0000_0000_0800_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 156-1 ; //100

      256'h0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 157-1 ; //99

      256'h0000_0000_0000_0000_0000_0000_2000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 158-1 ; //98

      256'h0000_0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 159-1 ; //97

      256'h0000_0000_0000_0000_0000_0000_8000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 160-1 ; //96

      256'h0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 161-1 ; //95

      256'h0000_0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 162-1 ; //94

      256'h0000_0000_0000_0000_0000_0004_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 163-1 ; //93

      256'h0000_0000_0000_0000_0000_0008_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 164-1 ; //92

      256'h0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 165-1 ; //91

      256'h0000_0000_0000_0000_0000_0020_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 166-1 ; //90

      256'h0000_0000_0000_0000_0000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 167-1 ; //89

      256'h0000_0000_0000_0000_0000_0080_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 168-1 ; //88

      256'h0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 169-1 ; //87

      256'h0000_0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 170-1 ; //86

      256'h0000_0000_0000_0000_0000_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 171-1 ; //85

      256'h0000_0000_0000_0000_0000_0800_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 172-1 ; //84

      256'h0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 173-1 ; //83

      256'h0000_0000_0000_0000_0000_2000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 174-1 ; //82

      256'h0000_0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 175-1 ; //81

      256'h0000_0000_0000_0000_0000_8000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 176-1 ; //80

      256'h0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 177-1 ; //79

      256'h0000_0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 178-1 ; //78

      256'h0000_0000_0000_0000_0004_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 179-1 ; //77

      256'h0000_0000_0000_0000_0008_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 180-1 ; //76

      256'h0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 181-1 ; //75

      256'h0000_0000_0000_0000_0020_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 182-1 ; //74

      256'h0000_0000_0000_0000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 183-1 ; //73

      256'h0000_0000_0000_0000_0080_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 184-1 ; //72

      256'h0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 185-1 ; //71

      256'h0000_0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 186-1 ; //70

      256'h0000_0000_0000_0000_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 187-1 ; //69

      256'h0000_0000_0000_0000_0800_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 188-1 ; //68

      256'h0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 189-1 ; //67

      256'h0000_0000_0000_0000_2000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 190-1 ; //66

      256'h0000_0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 191-1 ; //65

      256'h0000_0000_0000_0000_8000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 192-1 ; //64

      256'h0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 193-1 ; //63

      256'h0000_0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 194-1 ; //62

      256'h0000_0000_0000_0004_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 195-1 ; //61

      256'h0000_0000_0000_0008_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 196-1 ; //60

      256'h0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 197-1 ; //59

      256'h0000_0000_0000_0020_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 198-1 ; //58

      256'h0000_0000_0000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 199-1 ; //57

      256'h0000_0000_0000_0080_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 200-1 ; //56

      256'h0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 201-1 ; //55

      256'h0000_0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 202-1 ; //54

      256'h0000_0000_0000_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 203-1 ; //53

      256'h0000_0000_0000_0800_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 204-1 ; //52

      256'h0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 205-1 ; //51

      256'h0000_0000_0000_2000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 206-1 ; //50

      256'h0000_0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 207-1 ; //49

      256'h0000_0000_0000_8000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 208-1 ; //48

      256'h0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 209-1 ; //47

      256'h0000_0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 210-1 ; //46

      256'h0000_0000_0004_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 211-1 ; //45

      256'h0000_0000_0008_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 212-1 ; //44

      256'h0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 213-1 ; //43

      256'h0000_0000_0020_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 214-1 ; //42

      256'h0000_0000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 215-1 ; //41

      256'h0000_0000_0080_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 216-1 ; //40

      256'h0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 217-1 ; //39

      256'h0000_0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 218-1 ; //38

      256'h0000_0000_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 219-1 ; //37

      256'h0000_0000_0800_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 220-1 ; //36

      256'h0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 221-1 ; //35

      256'h0000_0000_2000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 222-1 ; //34

      256'h0000_0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 223-1 ; //33

      256'h0000_0000_8000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 224-1 ; //32

      256'h0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 225-1 ; //31

      256'h0000_0002_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 226-1 ; //30

      256'h0000_0004_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 227-1 ; //29

      256'h0000_0008_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 228-1 ; //28

      256'h0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 229-1 ; //27

      256'h0000_0020_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 230-1 ; //26

      256'h0000_0040_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 231-1 ; //25

      256'h0000_0080_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 232-1 ; //24

      256'h0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 233-1 ; //23

      256'h0000_0200_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 234-1 ; //22

      256'h0000_0400_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 235-1 ; //21

      256'h0000_0800_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 236-1 ; //20

      256'h0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 237-1 ; //19

      256'h0000_2000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 238-1 ; //18

      256'h0000_4000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 239-1 ; //17

      256'h0000_8000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 240-1 ; //16

      // 256'h0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: sel_enc = BASE + 242-1 ; //7

      default: sel_enc = BASE + 255;

    endcase
  end

endmodule : encoder_256_8
         
