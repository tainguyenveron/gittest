`include "sequence_read.sv"
`include "sequence_write.sv"
